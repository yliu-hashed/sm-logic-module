`default_nettype none

module top (
  input  [6:0] byte_i,
  (* color = "black" *)
  output reg [34:0] disp_o
  );

  /* ASCII TABLE -------------------------- */
  /*                                        */
  /*     0 1 2 3 4 5 6 7 8 9 A B C D E F    */
  /*  0                                     */
  /*  1                                     */
  /*  2    ! " # $ % & ' ( ) * + , - . /    */
  /*  3  0 1 2 3 4 5 6 7 8 9 : ; < = > ?    */
  /*  4  @ A B C D E F G H I J K L M N O    */
  /*  5  P Q R S T U V W X Y Z [ \ ] ^ _    */
  /*  6  ` a b c d e f g h i j k l m n o    */
  /*  8  p q r s t u v w x y z { | } ~      */
  /*                                        */
  /* -------------------------------------- */

  always @(byte_i) begin
    case (byte_i)
      default: disp_o <= {35{1'bX}}; // other characters are don't care
      7'h09: disp_o <= 35'h0; // horizontal tab
      7'h0B: disp_o <= 35'h0; // vertical tab
      7'h20: disp_o <= 35'h0; // spacebar
      // -----------------------------------------------------------------------
      // Specials
      // -----------------------------------------------------------------------
      7'h21: disp_o = { 5'b00100, // [!]
                        5'b00100,
                        5'b00100,
                        5'b00100,
                        5'b00100,
                        5'b00000,
                        5'b00100 };
      7'h22: disp_o = { 5'b01010, // ["]
                        5'b01010,
                        5'b00000,
                        5'b00000,
                        5'b00000,
                        5'b00000,
                        5'b00000 };
      7'h23: disp_o = { 5'b01010, // [#]
                        5'b01010,
                        5'b11111,
                        5'b01010,
                        5'b11111,
                        5'b01010,
                        5'b01010 };
      7'h24: disp_o = { 5'b00100, // [$]
                        5'b11111,
                        5'b10100,
                        5'b11111,
                        5'b00101,
                        5'b11111,
                        5'b00100 };
      7'h25: disp_o = { 5'b11001, // [%]
                        5'b11001,
                        5'b00010,
                        5'b00100,
                        5'b01000,
                        5'b10011,
                        5'b10011 };
      7'h26: disp_o = { 5'b01110, // [&]
                        5'b01010,
                        5'b00100,
                        5'b01101,
                        5'b10011,
                        5'b10001,
                        5'b01110 };
      7'h27: disp_o = { 5'b00100, // [']
                        5'b00100,
                        5'b00000,
                        5'b00000,
                        5'b00000,
                        5'b00000,
                        5'b00000 };
      7'h28: disp_o = { 5'b00010, // [(]
                        5'b00100,
                        5'b01000,
                        5'b01000,
                        5'b01000,
                        5'b00100,
                        5'b00010 };
      7'h29: disp_o = { 5'b01000, // [)]
                        5'b00100,
                        5'b00010,
                        5'b00010,
                        5'b00010,
                        5'b00100,
                        5'b01000 };
      7'h2A: disp_o = { 5'b00000, // [*]
                        5'b00100,
                        5'b10101,
                        5'b01110,
                        5'b10101,
                        5'b00100,
                        5'b00000 };
      7'h2B: disp_o = { 5'b00000, // [+]
                        5'b00100,
                        5'b00100,
                        5'b11111,
                        5'b00100,
                        5'b00100,
                        5'b00000 };
      7'h2C: disp_o = { 5'b00000, // [,]
                        5'b00000,
                        5'b00000,
                        5'b00000,
                        5'b00100,
                        5'b00100,
                        5'b01000 };
      7'h2D: disp_o = { 5'b00000, // [-]
                        5'b00000,
                        5'b00000,
                        5'b11111,
                        5'b00000,
                        5'b00000,
                        5'b00000 };
      7'h2E: disp_o = { 5'b00000, // [.]
                        5'b00000,
                        5'b00000,
                        5'b00000,
                        5'b00000,
                        5'b00000,
                        5'b00100 };
      7'h2F: disp_o = { 5'b00010, // [/]
                        5'b00010,
                        5'b00100,
                        5'b00100,
                        5'b00100,
                        5'b01000,
                        5'b01000 };
      // -----------------------------------------------------------------------
      // Numerical Digits
      // -----------------------------------------------------------------------
      7'h30: disp_o = { 5'b01110, // [0]
                        5'b10001,
                        5'b10011,
                        5'b10101,
                        5'b11001,
                        5'b10001,
                        5'b01110 };
      7'h31: disp_o = { 5'b00100, // [1]
                        5'b01100,
                        5'b00100,
                        5'b00100,
                        5'b00100,
                        5'b00100,
                        5'b11111 };
      7'h32: disp_o = { 5'b01110, // [2]
                        5'b10001,
                        5'b00001,
                        5'b00010,
                        5'b00100,
                        5'b01000,
                        5'b11111 };
      7'h33: disp_o = { 5'b01110, // [3]
                        5'b10001,
                        5'b00001,
                        5'b00110,
                        5'b00001,
                        5'b10001,
                        5'b01110 };
      7'h34: disp_o = { 5'b00010, // [4]
                        5'b00110,
                        5'b01010,
                        5'b10010,
                        5'b11111,
                        5'b00010,
                        5'b00010 };
      7'h35: disp_o = { 5'b11111, // [5]
                        5'b10000,
                        5'b11110,
                        5'b00001,
                        5'b00001,
                        5'b10001,
                        5'b01110 };
      7'h36: disp_o = { 5'b01110, // [6]
                        5'b10001,
                        5'b10000,
                        5'b11110,
                        5'b10001,
                        5'b10001,
                        5'b01110 };
      7'h37: disp_o = { 5'b11111, // [7]
                        5'b00001,
                        5'b00001,
                        5'b00010,
                        5'b00010,
                        5'b00100,
                        5'b00100 };
      7'h38: disp_o = { 5'b01110, // [8]
                        5'b10001,
                        5'b10001,
                        5'b01110,
                        5'b10001,
                        5'b10001,
                        5'b01110 };
      7'h39: disp_o = { 5'b01110, // [9]
                        5'b10001,
                        5'b10001,
                        5'b01111,
                        5'b00001,
                        5'b00010,
                        5'b01100 };
      // -----------------------------------------------------------------------
      // Specials After Numerical Digits
      // -----------------------------------------------------------------------
      7'h3A: disp_o = { 5'b00000, // [:]
                        5'b00000,
                        5'b00100,
                        5'b00000,
                        5'b00100,
                        5'b00000,
                        5'b00000 };
      7'h3B: disp_o = { 5'b00000, // [;]
                        5'b00000,
                        5'b00100,
                        5'b00000,
                        5'b00100,
                        5'b00100,
                        5'b01000 };
      7'h3C: disp_o = { 5'b00000, // [<]
                        5'b00010,
                        5'b00100,
                        5'b01000,
                        5'b00100,
                        5'b00010,
                        5'b00000 };
      7'h3D: disp_o = { 5'b00000, // [=]
                        5'b00000,
                        5'b01110,
                        5'b00000,
                        5'b01110,
                        5'b00000,
                        5'b00000 };
      7'h3E: disp_o = { 5'b00000, // [>]
                        5'b01000,
                        5'b00100,
                        5'b00010,
                        5'b00100,
                        5'b01000,
                        5'b00000 };
      7'h3F: disp_o = { 5'b01110, // [?]
                        5'b10001,
                        5'b00001,
                        5'b00010,
                        5'b00100,
                        5'b00000,
                        5'b00100 };
      7'h40: disp_o = { 5'b01110, // [@]
                        5'b10001,
                        5'b10111,
                        5'b10101,
                        5'b10111,
                        5'b10000,
                        5'b01110 };
      // -----------------------------------------------------------------------
      // Upper Cased Letters
      // -----------------------------------------------------------------------
      7'h41: disp_o = { 5'b01110, // [A]
                        5'b10001,
                        5'b10001,
                        5'b11111,
                        5'b10001,
                        5'b10001,
                        5'b10001 };
      7'h42: disp_o = { 5'b11110, // [B]
                        5'b10001,
                        5'b10001,
                        5'b11110,
                        5'b10001,
                        5'b10001,
                        5'b11110 };
      7'h43: disp_o = { 5'b01110, // [C]
                        5'b10001,
                        5'b10000,
                        5'b10000,
                        5'b10000,
                        5'b10001,
                        5'b01110 };
      7'h44: disp_o = { 5'b11110, // [D]
                        5'b10001,
                        5'b10001,
                        5'b10001,
                        5'b10001,
                        5'b10001,
                        5'b11110 };
      7'h45: disp_o = { 5'b11111, // [E]
                        5'b10000,
                        5'b10000,
                        5'b11110,
                        5'b10000,
                        5'b10000,
                        5'b11111 };
      7'h46: disp_o = { 5'b11111, // [F]
                        5'b10000,
                        5'b10000,
                        5'b11110,
                        5'b10000,
                        5'b10000,
                        5'b10000 };
      7'h47: disp_o = { 5'b01110, // [G]
                        5'b10001,
                        5'b10000,
                        5'b10011,
                        5'b10001,
                        5'b10001,
                        5'b01110 };
      7'h48: disp_o = { 5'b10001, // [H]
                        5'b10001,
                        5'b10001,
                        5'b11111,
                        5'b10001,
                        5'b10001,
                        5'b10001 };
      7'h49: disp_o = { 5'b01110, // [I]
                        5'b00100,
                        5'b00100,
                        5'b00100,
                        5'b00100,
                        5'b00100,
                        5'b01110 };
      7'h4A: disp_o = { 5'b01110, // [J]
                        5'b00010,
                        5'b00010,
                        5'b00010,
                        5'b10010,
                        5'b10010,
                        5'b01100 };
      7'h4B: disp_o = { 5'b10001, // [K]
                        5'b10001,
                        5'b10010,
                        5'b11100,
                        5'b10010,
                        5'b10001,
                        5'b10001 };
      7'h4C: disp_o = { 5'b10000, // [L]
                        5'b10000,
                        5'b10000,
                        5'b10000,
                        5'b10000,
                        5'b10000,
                        5'b11111 };
      7'h4D: disp_o = { 5'b10001, // [M]
                        5'b11011,
                        5'b10101,
                        5'b10001,
                        5'b10001,
                        5'b10001,
                        5'b10001 };
      7'h4E: disp_o = { 5'b10001, // [N]
                        5'b11001,
                        5'b10101,
                        5'b10011,
                        5'b10001,
                        5'b10001,
                        5'b10001 };
      7'h4F: disp_o = { 5'b01110, // [O]
                        5'b10001,
                        5'b10001,
                        5'b10001,
                        5'b10001,
                        5'b10001,
                        5'b01110 };
      7'h50: disp_o = { 5'b11110, // [P]
                        5'b10001,
                        5'b10001,
                        5'b11110,
                        5'b10000,
                        5'b10000,
                        5'b10000 };
      7'h51: disp_o = { 5'b01110, // [Q]
                        5'b10001,
                        5'b10001,
                        5'b10001,
                        5'b10101,
                        5'b10010,
                        5'b01101 };
      7'h52: disp_o = { 5'b01110, // [R]
                        5'b10001,
                        5'b10001,
                        5'b11110,
                        5'b10100,
                        5'b10010,
                        5'b10001 };
      7'h53: disp_o = { 5'b01110, // [S]
                        5'b10001,
                        5'b10000,
                        5'b01110,
                        5'b00001,
                        5'b10001,
                        5'b01110 };
      7'h54: disp_o = { 5'b11111, // [T]
                        5'b00100,
                        5'b00100,
                        5'b00100,
                        5'b00100,
                        5'b00100,
                        5'b00100 };
      7'h55: disp_o = { 5'b10001, // [U]
                        5'b10001,
                        5'b10001,
                        5'b10001,
                        5'b10001,
                        5'b10001,
                        5'b01110 };
      7'h56: disp_o = { 5'b10001, // [V]
                        5'b10001,
                        5'b10001,
                        5'b10001,
                        5'b01010,
                        5'b01010,
                        5'b00100 };
      7'h57: disp_o = { 5'b10001, // [W]
                        5'b10001,
                        5'b10001,
                        5'b10001,
                        5'b10101,
                        5'b10101,
                        5'b01010 };
      7'h58: disp_o = { 5'b10001, // [X]
                        5'b10001,
                        5'b01010,
                        5'b00100,
                        5'b01010,
                        5'b10001,
                        5'b10001 };
      7'h59: disp_o = { 5'b10001, // [Y]
                        5'b10001,
                        5'b01010,
                        5'b00100,
                        5'b00100,
                        5'b00100,
                        5'b00100 };
      7'h5A: disp_o = { 5'b11111, // [Z]
                        5'b00001,
                        5'b00010,
                        5'b00100,
                        5'b01000,
                        5'b10000,
                        5'b11111 };
      // -----------------------------------------------------------------------
      // Specials After Upper Cased Letters
      // -----------------------------------------------------------------------
      7'h5B: disp_o = { 5'b01110, // [[]
                        5'b01000,
                        5'b01000,
                        5'b01000,
                        5'b01000,
                        5'b01000,
                        5'b01110 };
      7'h5C: disp_o = { 5'b01000, // [\]
                        5'b01000,
                        5'b00100,
                        5'b00100,
                        5'b00100,
                        5'b00010,
                        5'b00010 };
      7'h5D: disp_o = { 5'b01110, // []]
                        5'b00010,
                        5'b00010,
                        5'b00010,
                        5'b00010,
                        5'b00010,
                        5'b01110 };
      7'h5E: disp_o = { 5'b00100, // [^]
                        5'b01010,
                        5'b00000,
                        5'b00000,
                        5'b00000,
                        5'b00000,
                        5'b00000 };
      7'h5F: disp_o = { 5'b00000, // [_]
                        5'b00000,
                        5'b00000,
                        5'b00000,
                        5'b00000,
                        5'b00000,
                        5'b11111 };
      7'h60: disp_o = { 5'b01000, // [`]
                        5'b00100,
                        5'b00000,
                        5'b00000,
                        5'b00000,
                        5'b00000,
                        5'b00000 };
      // -----------------------------------------------------------------------
      // Lower Cased Letters
      // -----------------------------------------------------------------------
      7'h61: disp_o = { 5'b00000, // [a]
                        5'b00000,
                        5'b01110,
                        5'b00001,
                        5'b01111,
                        5'b10001,
                        5'b01110 };
      7'h62: disp_o = { 5'b10000, // [b]
                        5'b10000,
                        5'b11110,
                        5'b10001,
                        5'b10001,
                        5'b10001,
                        5'b11110 };
      7'h63: disp_o = { 5'b00000, // [c]
                        5'b00000,
                        5'b01111,
                        5'b10000,
                        5'b10000,
                        5'b10000,
                        5'b01111 };
      7'h64: disp_o = { 5'b00001, // [d]
                        5'b00001,
                        5'b01111,
                        5'b10001,
                        5'b10001,
                        5'b10001,
                        5'b01111 };
      7'h65: disp_o = { 5'b00000, // [e]
                        5'b00000,
                        5'b01110,
                        5'b10001,
                        5'b11110,
                        5'b10000,
                        5'b01110 };
      7'h66: disp_o = { 5'b00110, // [f]
                        5'b01000,
                        5'b11111,
                        5'b01000,
                        5'b01000,
                        5'b01000,
                        5'b01000 };
      7'h67: disp_o = { 5'b00000, // [g]
                        5'b00000,
                        5'b01110,
                        5'b10001,
                        5'b01111,
                        5'b00001,
                        5'b01110 };
      7'h68: disp_o = { 5'b10000, // [h]
                        5'b10000,
                        5'b11110,
                        5'b10001,
                        5'b10001,
                        5'b10001,
                        5'b10001 };
      7'h69: disp_o = { 5'b00100, // [i]
                        5'b00000,
                        5'b11100,
                        5'b00100,
                        5'b00100,
                        5'b00100,
                        5'b11111 };
      7'h6A: disp_o = { 5'b00010, // [j]
                        5'b00000,
                        5'b01110,
                        5'b00010,
                        5'b00010,
                        5'b10010,
                        5'b01100 };
      7'h6B: disp_o = { 5'b10000, // [k]
                        5'b10000,
                        5'b10010,
                        5'b11100,
                        5'b10010,
                        5'b10001,
                        5'b10001 };
      7'h6C: disp_o = { 5'b11100, // [l]
                        5'b00100,
                        5'b00100,
                        5'b00100,
                        5'b00100,
                        5'b00100,
                        5'b00011 };
      7'h6D: disp_o = { 5'b00000, // [m]
                        5'b00000,
                        5'b01010,
                        5'b10101,
                        5'b10101,
                        5'b10101,
                        5'b10101 };
      7'h6E: disp_o = { 5'b00000, // [n]
                        5'b00000,
                        5'b11110,
                        5'b10001,
                        5'b10001,
                        5'b10001,
                        5'b10001 };
      7'h6F: disp_o = { 5'b00000, // [o]
                        5'b00000,
                        5'b01110,
                        5'b10001,
                        5'b10001,
                        5'b10001,
                        5'b01110 };
      7'h70: disp_o = { 5'b00000, // [p]
                        5'b00000,
                        5'b11110,
                        5'b10001,
                        5'b11110,
                        5'b10000,
                        5'b10000 };
      7'h71: disp_o = { 5'b00000, // [q]
                        5'b00000,
                        5'b01111,
                        5'b10001,
                        5'b01111,
                        5'b00001,
                        5'b00001 };
      7'h72: disp_o = { 5'b00000, // [r]
                        5'b00000,
                        5'b10110,
                        5'b11001,
                        5'b10000,
                        5'b10000,
                        5'b10000 };
      7'h73: disp_o = { 5'b00000, // [s]
                        5'b00000,
                        5'b01110,
                        5'b10000,
                        5'b01110,
                        5'b00001,
                        5'b01110 };
      7'h74: disp_o = { 5'b01000, // [t]
                        5'b01000,
                        5'b11111,
                        5'b01000,
                        5'b01000,
                        5'b01000,
                        5'b00111 };
      7'h75: disp_o = { 5'b00000, // [u]
                        5'b00000,
                        5'b10001,
                        5'b10001,
                        5'b10001,
                        5'b10001,
                        5'b01110 };
      7'h76: disp_o = { 5'b00000, // [v]
                        5'b00000,
                        5'b10001,
                        5'b10001,
                        5'b01010,
                        5'b01010,
                        5'b00100 };
      7'h77: disp_o = { 5'b00000, // [w]
                        5'b00000,
                        5'b10001,
                        5'b10001,
                        5'b10101,
                        5'b10101,
                        5'b01010 };
      7'h78: disp_o = { 5'b00000, // [x]
                        5'b00000,
                        5'b10001,
                        5'b01010,
                        5'b00100,
                        5'b01010,
                        5'b10001 };
      7'h79: disp_o = { 5'b00000, // [y]
                        5'b00000,
                        5'b10001,
                        5'b10001,
                        5'b01111,
                        5'b00001,
                        5'b01110 };
      7'h7A: disp_o = { 5'b00000, // [z]
                        5'b00000,
                        5'b11111,
                        5'b00010,
                        5'b00100,
                        5'b01000,
                        5'b11111 };
      // -----------------------------------------------------------------------
      // Specials After Lower Cased Letters
      // -----------------------------------------------------------------------
      7'h7B: disp_o = { 5'b00010, // [{]
                        5'b00100,
                        5'b00100,
                        5'b01000,
                        5'b00100,
                        5'b00100,
                        5'b00010 };
      7'h7C: disp_o = { 5'b00100, // [|]
                        5'b00100,
                        5'b00100,
                        5'b00100,
                        5'b00100,
                        5'b00100,
                        5'b00100 };
      7'h7D: disp_o = { 5'b01000, // [}]
                        5'b00100,
                        5'b00100,
                        5'b00010,
                        5'b00100,
                        5'b00100,
                        5'b01000 };
      7'h7E: disp_o = { 5'b00000, // [~]
                        5'b00000,
                        5'b01000,
                        5'b10101,
                        5'b00010,
                        5'b00000,
                        5'b00000 };
    endcase
  end
endmodule
